*Micro-Cap Tube Library
*http://www.spectrum-soft.com


*Beam Power Tetrode
*Based on the Norman Koren model with IG2 adaptation from Alexander Gurskii
.SUBCKT 4X150 1 2 3 4 ; P G1 C G2
+ PARAMS: MU=40.881 EX=645.155m KG1=20.02 KG2=437.262 KP=27.399 KVB=58.685
+ CCG=16P CPG1=.03P CCP=4.4P RGI=2K
RE1 7 0 1G
RE2 8 3 1G
E1 7 0 VALUE={V(4,3)/KP*LN(1+EXP((1/MU+V(2,3)/V(4,3))*KP))}
G1 1 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG1*ATAN(V(1,3)/KVB)}
G2 8 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG2*(2.5708-ATAN(V(1,3)/KVB))}
E2 8 4 VALUE={0}
RCP 1 3 1G
C1 2 3 {CCG} ; CATHODE-GRID 1 Capacitance
C2 1 2 {CPG1} ; GRID 1-PLATE Capacitance
C3 1 3 {CCP} ; CATHODE-PLATE Capacitance
R1 2 5 {RGI} ; FOR GRID CURRENT
D3 5 3 DX ; FOR GRID CURRENT
.MODEL DX D(IS=1N RS=1 CJO=10PF TT=1N)
.ENDS

*High Performance Audio Beam Power Tetrode
*Based on the Norman Koren model with IG2 adaptation from Alexander Gurskii
.SUBCKT 6L6GC 1 2 3 4 ; P G1 C G2
+ PARAMS: MU=19.684 EX=1.519 KG1=1.15K KG2=3000 KP=18.899 KVB=13.847
+ CCG=10P CPG1=.6P CCP=6.5P RGI=2K
RE1 7 0 1G
RE2 8 3 1G
E1 7 0 VALUE={V(4,3)/KP*LN(1+EXP((1/MU+V(2,3)/V(4,3))*KP))}
G1 1 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG1*ATAN(V(1,3)/KVB)}
G2 8 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG2*(2.5708-ATAN(V(1,3)/KVB))}
E2 8 4 VALUE={0}
RCP 1 3 1G ; FOR CONVERGENCE
C1 2 3 {CCG} ; CATHODE-GRID 1
C2 1 2 {CPG1} ; GRID 1-PLATE
C3 1 3 {CCP} ; CATHODE-PLATE
R1 2 5 {RGI} ; FOR GRID CURRENT
D3 5 3 DX ; FOR GRID CURRENT
.MODEL DX D(IS=1N RS=1 CJO=10PF TT=1N)
.ENDS

*High Performance Audio Power Pentode
*Based on the Norman Koren model with IG2 adaptation from Alexander Gurskii
.SUBCKT EL34 1 2 3 4 ; P G1 C G2
+ PARAMS: MU=9.67 EX=1.63 KG1=2.109K KG2=4100 KP=70.931 KVB=26.643
+ CCG=15.2P CPG1=1.1P CCP=8.4P RGI=2K
RE1 7 0 1G
RE2 8 3 1G
E1 7 0 VALUE={V(4,3)/KP*LN(1+EXP((1/MU+V(2,3)/V(4,3))*KP))}
G1 1 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG1*ATAN(V(1,3)/KVB)}
G2 8 3 VALUE={(PWR(V(7),EX)+PWRS(V(7),EX))/KG2*(2.5708-ATAN(V(1,3)/KVB))}
E2 8 4 VALUE={0}
RCP 1 3 1G ; FOR CONVERGENCE
C1 2 3 {CCG} ; CATHODE-GRID 1
C2 1 2 {CPG1} ; GRID 1-PLATE
C3 1 3 {CCP} ; CATHODE-PLATE
R1 2 5 {RGI} ; FOR GRID CURRENT
D3 5 3 DX ; FOR GRID CURRENT
.MODEL DX D(IS=1N RS=1 CJO=10PF TT=1N)
.ENDS
